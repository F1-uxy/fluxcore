module cpu (
    input logic clk,
    input logic reset,
    output logic [7:0] addr_bus,
    inout
);
    
endmodule